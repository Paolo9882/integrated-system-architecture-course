library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Dadda Tree
entity dadda_tree is
	port(
		pp0: in std_logic_vector(36 downto 0); --partial products
		pp1: in std_logic_vector(36 downto 0);
		pp2: in std_logic_vector(36 downto 0);
		pp3: in std_logic_vector(36 downto 0);
		pp4: in std_logic_vector(36 downto 0);
		pp5: in std_logic_vector(36 downto 0);
		pp6: in std_logic_vector(36 downto 0);
		pp7: in std_logic_vector(36 downto 0);
		pp8: in std_logic_vector(36 downto 0);
		pp9: in std_logic_vector(36 downto 0);
		pp10: in std_logic_vector(36 downto 0);
		pp11: in std_logic_vector(36 downto 0);
		pp12: in std_logic_vector(36 downto 0);
		pp13: in std_logic_vector(36 downto 0);
		pp14: in std_logic_vector(36 downto 0);
		pp15: in std_logic_vector(36 downto 0);
		pp16: in std_logic_vector(36 downto 0);		
		final0: out std_logic_vector(63 downto 0); --final two addends
		final1: out std_logic_vector(63 downto 0)
	);
end dadda_tree;

architecture structural of dadda_tree is

	--partial signals and port map described by dadda_tree_generator.py
	signal pp17	: std_logic_vector(63 downto 0);
	signal pp18	: std_logic_vector(63 downto 0);
	signal pp19	: std_logic_vector(63 downto 0);
	signal pp20	: std_logic_vector(63 downto 0);
	signal pp21	: std_logic_vector(63 downto 0);
	signal pp22	: std_logic_vector(63 downto 0);
	signal pp23	: std_logic_vector(63 downto 0);
	signal pp24	: std_logic_vector(63 downto 0);
	signal pp25	: std_logic_vector(63 downto 0);
	signal pp26	: std_logic_vector(63 downto 0);
	signal pp27	: std_logic_vector(63 downto 0);
	signal pp28	: std_logic_vector(63 downto 0);
	signal pp29	: std_logic_vector(63 downto 0);
	signal pp30	: std_logic_vector(63 downto 0);
	signal pp31	: std_logic_vector(63 downto 0);
	signal pp32	: std_logic_vector(63 downto 0);
	signal pp33	: std_logic_vector(63 downto 0);
	signal pp34	: std_logic_vector(63 downto 0);
	signal pp35	: std_logic_vector(63 downto 0);
	signal pp36	: std_logic_vector(63 downto 0);
	signal pp37	: std_logic_vector(63 downto 0);
	signal pp38	: std_logic_vector(63 downto 0);
	signal pp39	: std_logic_vector(63 downto 0);
	signal pp40	: std_logic_vector(63 downto 0);
	signal pp41	: std_logic_vector(63 downto 0);
	signal pp42	: std_logic_vector(63 downto 0);
	signal pp43	: std_logic_vector(63 downto 0);
	signal pp44	: std_logic_vector(63 downto 0);
	signal pp45	: std_logic_vector(63 downto 0);
	signal pp46	: std_logic_vector(63 downto 0);

	--components declaration
	component half_adder is
		port(
			a, b : in std_logic; --addends
			s, cout : out std_logic --sum and carry out
		);
	end component;

	component full_adder is
		port(
			a, b, cin : in std_logic; --addends
			s, cout : out std_logic --sum and carry out
		);
	end component;

	begin

	HA0: half_adder port map(
		a => pp0(24),
		b => pp1(24),
		s => pp17(24),
		cout => pp17(25)
		);

	HA1: half_adder port map(
		a => pp0(25),
		b => pp1(25),
		s => pp18(25),
		cout => pp17(26)
		);

	FA0: full_adder port map(
		a => pp0(26),
		b => pp1(26),
		cin => pp2(24),
		s => pp18(26),
		cout => pp17(27)
		);

	HA2: half_adder port map(
		a => pp3(22),
		b => pp4(20),
		s => pp19(26),
		cout => pp18(27)
		);

	FA1: full_adder port map(
		a => pp0(27),
		b => pp1(27),
		cin => pp2(25),
		s => pp19(27),
		cout => pp17(28)
		);

	HA3: half_adder port map(
		a => pp3(23),
		b => pp4(21),
		s => pp20(27),
		cout => pp18(28)
		);

	FA2: full_adder port map(
		a => pp0(28),
		b => pp1(28),
		cin => pp2(26),
		s => pp19(28),
		cout => pp17(29)
		);

	FA3: full_adder port map(
		a => pp3(24),
		b => pp4(22),
		cin => pp5(20),
		s => pp20(28),
		cout => pp18(29)
		);

	HA4: half_adder port map(
		a => pp6(18),
		b => pp7(16),
		s => pp21(28),
		cout => pp19(29)
		);

	FA4: full_adder port map(
		a => pp0(29),
		b => pp1(29),
		cin => pp2(27),
		s => pp20(29),
		cout => pp17(30)
		);

	FA5: full_adder port map(
		a => pp3(25),
		b => pp4(23),
		cin => pp5(21),
		s => pp21(29),
		cout => pp18(30)
		);

	HA5: half_adder port map(
		a => pp6(19),
		b => pp7(17),
		s => pp22(29),
		cout => pp19(30)
		);

	FA6: full_adder port map(
		a => pp0(30),
		b => pp1(30),
		cin => pp2(28),
		s => pp20(30),
		cout => pp17(31)
		);

	FA7: full_adder port map(
		a => pp3(26),
		b => pp4(24),
		cin => pp5(22),
		s => pp21(30),
		cout => pp18(31)
		);

	FA8: full_adder port map(
		a => pp6(20),
		b => pp7(18),
		cin => pp8(16),
		s => pp22(30),
		cout => pp19(31)
		);

	HA6: half_adder port map(
		a => pp9(14),
		b => pp10(12),
		s => pp23(30),
		cout => pp20(31)
		);

	FA9: full_adder port map(
		a => pp0(31),
		b => pp1(31),
		cin => pp2(29),
		s => pp21(31),
		cout => pp17(32)
		);

	FA10: full_adder port map(
		a => pp3(27),
		b => pp4(25),
		cin => pp5(23),
		s => pp22(31),
		cout => pp18(32)
		);

	FA11: full_adder port map(
		a => pp6(21),
		b => pp7(19),
		cin => pp8(17),
		s => pp23(31),
		cout => pp19(32)
		);

	HA7: half_adder port map(
		a => pp9(15),
		b => pp10(13),
		s => pp24(31),
		cout => pp20(32)
		);

	FA12: full_adder port map(
		a => pp0(32),
		b => pp1(32),
		cin => pp2(30),
		s => pp21(32),
		cout => pp17(33)
		);

	FA13: full_adder port map(
		a => pp3(28),
		b => pp4(26),
		cin => pp5(24),
		s => pp22(32),
		cout => pp18(33)
		);

	FA14: full_adder port map(
		a => pp6(22),
		b => pp7(20),
		cin => pp8(18),
		s => pp23(32),
		cout => pp19(33)
		);

	FA15: full_adder port map(
		a => pp9(16),
		b => pp10(14),
		cin => pp11(12),
		s => pp24(32),
		cout => pp20(33)
		);

	FA16: full_adder port map(
		a => pp0(33),
		b => pp1(33),
		cin => pp2(31),
		s => pp21(33),
		cout => pp17(34)
		);

	FA17: full_adder port map(
		a => pp3(29),
		b => pp4(27),
		cin => pp5(25),
		s => pp22(33),
		cout => pp18(34)
		);

	FA18: full_adder port map(
		a => pp6(23),
		b => pp7(21),
		cin => pp8(19),
		s => pp23(33),
		cout => pp19(34)
		);

	FA19: full_adder port map(
		a => pp9(17),
		b => pp10(15),
		cin => pp11(13),
		s => pp24(33),
		cout => pp20(34)
		);

	FA20: full_adder port map(
		a => pp0(34),
		b => pp1(34),
		cin => pp2(32),
		s => pp21(34),
		cout => pp17(35)
		);

	FA21: full_adder port map(
		a => pp3(30),
		b => pp4(28),
		cin => pp5(26),
		s => pp22(34),
		cout => pp18(35)
		);

	FA22: full_adder port map(
		a => pp6(24),
		b => pp7(22),
		cin => pp8(20),
		s => pp23(34),
		cout => pp19(35)
		);

	FA23: full_adder port map(
		a => pp9(18),
		b => pp10(16),
		cin => pp11(14),
		s => pp24(34),
		cout => pp20(35)
		);

	FA24: full_adder port map(
		a => pp0(35),
		b => pp1(35),
		cin => pp2(33),
		s => pp21(35),
		cout => pp17(36)
		);

	FA25: full_adder port map(
		a => pp3(31),
		b => pp4(29),
		cin => pp5(27),
		s => pp22(35),
		cout => pp18(36)
		);

	FA26: full_adder port map(
		a => pp6(25),
		b => pp7(23),
		cin => pp8(21),
		s => pp23(35),
		cout => pp19(36)
		);

	FA27: full_adder port map(
		a => pp9(19),
		b => pp10(17),
		cin => pp11(15),
		s => pp24(35),
		cout => pp20(36)
		);

	FA28: full_adder port map(
		a => pp1(36),
		b => pp2(34),
		cin => pp3(32),
		s => pp21(36),
		cout => pp17(37)
		);

	FA29: full_adder port map(
		a => pp4(30),
		b => pp5(28),
		cin => pp6(26),
		s => pp22(36),
		cout => pp18(37)
		);

	FA30: full_adder port map(
		a => pp7(24),
		b => pp8(22),
		cin => pp9(20),
		s => pp23(36),
		cout => pp19(37)
		);

	HA8: half_adder port map(
		a => pp10(18),
		b => pp11(16),
		s => pp24(36),
		cout => pp20(37)
		);

	FA31: full_adder port map(
		a => pp2(35),
		b => pp3(33),
		cin => pp4(31),
		s => pp21(37),
		cout => pp17(38)
		);

	FA32: full_adder port map(
		a => pp5(29),
		b => pp6(27),
		cin => pp7(25),
		s => pp22(37),
		cout => pp18(38)
		);

	FA33: full_adder port map(
		a => pp8(23),
		b => pp9(21),
		cin => pp10(19),
		s => pp23(37),
		cout => pp19(38)
		);

	FA34: full_adder port map(
		a => pp2(36),
		b => pp3(34),
		cin => pp4(32),
		s => pp20(38),
		cout => pp17(39)
		);

	FA35: full_adder port map(
		a => pp5(30),
		b => pp6(28),
		cin => pp7(26),
		s => pp21(38),
		cout => pp18(39)
		);

	HA9: half_adder port map(
		a => pp8(24),
		b => pp9(22),
		s => pp22(38),
		cout => pp19(39)
		);

	FA36: full_adder port map(
		a => pp3(35),
		b => pp4(33),
		cin => pp5(31),
		s => pp20(39),
		cout => pp17(40)
		);

	FA37: full_adder port map(
		a => pp6(29),
		b => pp7(27),
		cin => pp8(25),
		s => pp21(39),
		cout => pp18(40)
		);

	FA38: full_adder port map(
		a => pp3(36),
		b => pp4(34),
		cin => pp5(32),
		s => pp19(40),
		cout => pp17(41)
		);

	HA10: half_adder port map(
		a => pp6(30),
		b => pp7(28),
		s => pp20(40),
		cout => pp18(41)
		);

	FA39: full_adder port map(
		a => pp4(35),
		b => pp5(33),
		cin => pp6(31),
		s => pp19(41),
		cout => pp17(42)
		);

	HA11: half_adder port map(
		a => pp4(36),
		b => pp5(34),
		s => pp18(42),
		cout => pp17(43)
		);

	HA12: half_adder port map(
		a => pp0(16),
		b => pp1(16),
		s => pp25(16),
		cout => pp25(17)
		);

	HA13: half_adder port map(
		a => pp0(17),
		b => pp1(17),
		s => pp26(17),
		cout => pp25(18)
		);

	FA40: full_adder port map(
		a => pp0(18),
		b => pp1(18),
		cin => pp2(16),
		s => pp26(18),
		cout => pp25(19)
		);

	HA14: half_adder port map(
		a => pp3(14),
		b => pp4(12),
		s => pp27(18),
		cout => pp26(19)
		);

	FA41: full_adder port map(
		a => pp0(19),
		b => pp1(19),
		cin => pp2(17),
		s => pp27(19),
		cout => pp25(20)
		);

	HA15: half_adder port map(
		a => pp3(15),
		b => pp4(13),
		s => pp28(19),
		cout => pp26(20)
		);

	FA42: full_adder port map(
		a => pp0(20),
		b => pp1(20),
		cin => pp2(18),
		s => pp27(20),
		cout => pp25(21)
		);

	FA43: full_adder port map(
		a => pp3(16),
		b => pp4(14),
		cin => pp5(12),
		s => pp28(20),
		cout => pp26(21)
		);

	HA16: half_adder port map(
		a => pp6(10),
		b => pp7(8),
		s => pp29(20),
		cout => pp27(21)
		);

	FA44: full_adder port map(
		a => pp0(21),
		b => pp1(21),
		cin => pp2(19),
		s => pp28(21),
		cout => pp25(22)
		);

	FA45: full_adder port map(
		a => pp3(17),
		b => pp4(15),
		cin => pp5(13),
		s => pp29(21),
		cout => pp26(22)
		);

	HA17: half_adder port map(
		a => pp6(11),
		b => pp7(9),
		s => pp30(21),
		cout => pp27(22)
		);

	FA46: full_adder port map(
		a => pp0(22),
		b => pp1(22),
		cin => pp2(20),
		s => pp28(22),
		cout => pp25(23)
		);

	FA47: full_adder port map(
		a => pp3(18),
		b => pp4(16),
		cin => pp5(14),
		s => pp29(22),
		cout => pp26(23)
		);

	FA48: full_adder port map(
		a => pp6(12),
		b => pp7(10),
		cin => pp8(8),
		s => pp30(22),
		cout => pp27(23)
		);

	HA18: half_adder port map(
		a => pp9(6),
		b => pp10(4),
		s => pp31(22),
		cout => pp28(23)
		);

	FA49: full_adder port map(
		a => pp0(23),
		b => pp1(23),
		cin => pp2(21),
		s => pp29(23),
		cout => pp25(24)
		);

	FA50: full_adder port map(
		a => pp3(19),
		b => pp4(17),
		cin => pp5(15),
		s => pp30(23),
		cout => pp26(24)
		);

	FA51: full_adder port map(
		a => pp6(13),
		b => pp7(11),
		cin => pp8(9),
		s => pp31(23),
		cout => pp27(24)
		);

	HA19: half_adder port map(
		a => pp9(7),
		b => pp10(5),
		s => pp32(23),
		cout => pp28(24)
		);

	FA52: full_adder port map(
		a => pp2(22),
		b => pp3(20),
		cin => pp4(18),
		s => pp29(24),
		cout => pp25(25)
		);

	FA53: full_adder port map(
		a => pp5(16),
		b => pp6(14),
		cin => pp7(12),
		s => pp30(24),
		cout => pp26(25)
		);

	FA54: full_adder port map(
		a => pp8(10),
		b => pp9(8),
		cin => pp10(6),
		s => pp31(24),
		cout => pp27(25)
		);

	FA55: full_adder port map(
		a => pp11(4),
		b => pp12(2),
		cin => pp13(0),
		s => pp32(24),
		cout => pp28(25)
		);

	FA56: full_adder port map(
		a => pp2(23),
		b => pp3(21),
		cin => pp4(19),
		s => pp29(25),
		cout => pp25(26)
		);

	FA57: full_adder port map(
		a => pp5(17),
		b => pp6(15),
		cin => pp7(13),
		s => pp30(25),
		cout => pp26(26)
		);

	FA58: full_adder port map(
		a => pp8(11),
		b => pp9(9),
		cin => pp10(7),
		s => pp31(25),
		cout => pp27(26)
		);

	FA59: full_adder port map(
		a => pp11(5),
		b => pp12(3),
		cin => pp17(25),
		s => pp32(25),
		cout => pp28(26)
		);

	FA60: full_adder port map(
		a => pp5(18),
		b => pp6(16),
		cin => pp7(14),
		s => pp29(26),
		cout => pp25(27)
		);

	FA61: full_adder port map(
		a => pp8(12),
		b => pp9(10),
		cin => pp10(8),
		s => pp30(26),
		cout => pp26(27)
		);

	FA62: full_adder port map(
		a => pp11(6),
		b => pp12(4),
		cin => pp13(2),
		s => pp31(26),
		cout => pp27(27)
		);

	FA63: full_adder port map(
		a => pp14(0),
		b => pp17(26),
		cin => pp18(26),
		s => pp32(26),
		cout => pp28(27)
		);

	FA64: full_adder port map(
		a => pp5(19),
		b => pp6(17),
		cin => pp7(15),
		s => pp29(27),
		cout => pp25(28)
		);

	FA65: full_adder port map(
		a => pp8(13),
		b => pp9(11),
		cin => pp10(9),
		s => pp30(27),
		cout => pp26(28)
		);

	FA66: full_adder port map(
		a => pp11(7),
		b => pp12(5),
		cin => pp13(3),
		s => pp31(27),
		cout => pp27(28)
		);

	FA67: full_adder port map(
		a => pp17(27),
		b => pp18(27),
		cin => pp19(27),
		s => pp32(27),
		cout => pp28(28)
		);

	FA68: full_adder port map(
		a => pp8(14),
		b => pp9(12),
		cin => pp10(10),
		s => pp29(28),
		cout => pp25(29)
		);

	FA69: full_adder port map(
		a => pp11(8),
		b => pp12(6),
		cin => pp13(4),
		s => pp30(28),
		cout => pp26(29)
		);

	FA70: full_adder port map(
		a => pp14(2),
		b => pp15(0),
		cin => pp17(28),
		s => pp31(28),
		cout => pp27(29)
		);

	FA71: full_adder port map(
		a => pp18(28),
		b => pp19(28),
		cin => pp20(28),
		s => pp32(28),
		cout => pp28(29)
		);

	FA72: full_adder port map(
		a => pp8(15),
		b => pp9(13),
		cin => pp10(11),
		s => pp29(29),
		cout => pp25(30)
		);

	FA73: full_adder port map(
		a => pp11(9),
		b => pp12(7),
		cin => pp13(5),
		s => pp30(29),
		cout => pp26(30)
		);

	FA74: full_adder port map(
		a => pp14(3),
		b => pp17(29),
		cin => pp18(29),
		s => pp31(29),
		cout => pp27(30)
		);

	FA75: full_adder port map(
		a => pp19(29),
		b => pp20(29),
		cin => pp21(29),
		s => pp32(29),
		cout => pp28(30)
		);

	FA76: full_adder port map(
		a => pp11(10),
		b => pp12(8),
		cin => pp13(6),
		s => pp29(30),
		cout => pp25(31)
		);

	FA77: full_adder port map(
		a => pp14(4),
		b => pp15(2),
		cin => pp16(0),
		s => pp30(30),
		cout => pp26(31)
		);

	FA78: full_adder port map(
		a => pp17(30),
		b => pp18(30),
		cin => pp19(30),
		s => pp31(30),
		cout => pp27(31)
		);

	FA79: full_adder port map(
		a => pp20(30),
		b => pp21(30),
		cin => pp22(30),
		s => pp32(30),
		cout => pp28(31)
		);

	FA80: full_adder port map(
		a => pp11(11),
		b => pp12(9),
		cin => pp13(7),
		s => pp29(31),
		cout => pp25(32)
		);

	FA81: full_adder port map(
		a => pp14(5),
		b => pp15(3),
		cin => pp17(31),
		s => pp30(31),
		cout => pp26(32)
		);

	FA82: full_adder port map(
		a => pp18(31),
		b => pp19(31),
		cin => pp20(31),
		s => pp31(31),
		cout => pp27(32)
		);

	FA83: full_adder port map(
		a => pp21(31),
		b => pp22(31),
		cin => pp23(31),
		s => pp32(31),
		cout => pp28(32)
		);

	FA84: full_adder port map(
		a => pp12(10),
		b => pp13(8),
		cin => pp14(6),
		s => pp29(32),
		cout => pp25(33)
		);

	FA85: full_adder port map(
		a => pp15(4),
		b => pp16(2),
		cin => pp17(32),
		s => pp30(32),
		cout => pp26(33)
		);

	FA86: full_adder port map(
		a => pp18(32),
		b => pp19(32),
		cin => pp20(32),
		s => pp31(32),
		cout => pp27(33)
		);

	FA87: full_adder port map(
		a => pp21(32),
		b => pp22(32),
		cin => pp23(32),
		s => pp32(32),
		cout => pp28(33)
		);

	FA88: full_adder port map(
		a => pp12(11),
		b => pp13(9),
		cin => pp14(7),
		s => pp29(33),
		cout => pp25(34)
		);

	FA89: full_adder port map(
		a => pp15(5),
		b => pp16(3),
		cin => pp17(33),
		s => pp30(33),
		cout => pp26(34)
		);

	FA90: full_adder port map(
		a => pp18(33),
		b => pp19(33),
		cin => pp20(33),
		s => pp31(33),
		cout => pp27(34)
		);

	FA91: full_adder port map(
		a => pp21(33),
		b => pp22(33),
		cin => pp23(33),
		s => pp32(33),
		cout => pp28(34)
		);

	FA92: full_adder port map(
		a => pp12(12),
		b => pp13(10),
		cin => pp14(8),
		s => pp29(34),
		cout => pp25(35)
		);

	FA93: full_adder port map(
		a => pp15(6),
		b => pp16(4),
		cin => pp17(34),
		s => pp30(34),
		cout => pp26(35)
		);

	FA94: full_adder port map(
		a => pp18(34),
		b => pp19(34),
		cin => pp20(34),
		s => pp31(34),
		cout => pp27(35)
		);

	FA95: full_adder port map(
		a => pp21(34),
		b => pp22(34),
		cin => pp23(34),
		s => pp32(34),
		cout => pp28(35)
		);

	FA96: full_adder port map(
		a => pp12(13),
		b => pp13(11),
		cin => pp14(9),
		s => pp29(35),
		cout => pp25(36)
		);

	FA97: full_adder port map(
		a => pp15(7),
		b => pp16(5),
		cin => pp17(35),
		s => pp30(35),
		cout => pp26(36)
		);

	FA98: full_adder port map(
		a => pp18(35),
		b => pp19(35),
		cin => pp20(35),
		s => pp31(35),
		cout => pp27(36)
		);

	FA99: full_adder port map(
		a => pp21(35),
		b => pp22(35),
		cin => pp23(35),
		s => pp32(35),
		cout => pp28(36)
		);

	FA100: full_adder port map(
		a => pp12(14),
		b => pp13(12),
		cin => pp14(10),
		s => pp29(36),
		cout => pp25(37)
		);

	FA101: full_adder port map(
		a => pp15(8),
		b => pp16(6),
		cin => pp17(36),
		s => pp30(36),
		cout => pp26(37)
		);

	FA102: full_adder port map(
		a => pp18(36),
		b => pp19(36),
		cin => pp20(36),
		s => pp31(36),
		cout => pp27(37)
		);

	FA103: full_adder port map(
		a => pp21(36),
		b => pp22(36),
		cin => pp23(36),
		s => pp32(36),
		cout => pp28(37)
		);

	FA104: full_adder port map(
		a => pp11(17),
		b => pp12(15),
		cin => pp13(13),
		s => pp29(37),
		cout => pp25(38)
		);

	FA105: full_adder port map(
		a => pp14(11),
		b => pp15(9),
		cin => pp16(7),
		s => pp30(37),
		cout => pp26(38)
		);

	FA106: full_adder port map(
		a => pp17(37),
		b => pp18(37),
		cin => pp19(37),
		s => pp31(37),
		cout => pp27(38)
		);

	FA107: full_adder port map(
		a => pp20(37),
		b => pp21(37),
		cin => pp22(37),
		s => pp32(37),
		cout => pp28(38)
		);

	FA108: full_adder port map(
		a => pp10(20),
		b => pp11(18),
		cin => pp12(16),
		s => pp29(38),
		cout => pp25(39)
		);

	FA109: full_adder port map(
		a => pp13(14),
		b => pp14(12),
		cin => pp15(10),
		s => pp30(38),
		cout => pp26(39)
		);

	FA110: full_adder port map(
		a => pp16(8),
		b => pp17(38),
		cin => pp18(38),
		s => pp31(38),
		cout => pp27(39)
		);

	FA111: full_adder port map(
		a => pp19(38),
		b => pp20(38),
		cin => pp21(38),
		s => pp32(38),
		cout => pp28(39)
		);

	FA112: full_adder port map(
		a => pp9(23),
		b => pp10(21),
		cin => pp11(19),
		s => pp29(39),
		cout => pp25(40)
		);

	FA113: full_adder port map(
		a => pp12(17),
		b => pp13(15),
		cin => pp14(13),
		s => pp30(39),
		cout => pp26(40)
		);

	FA114: full_adder port map(
		a => pp15(11),
		b => pp16(9),
		cin => pp17(39),
		s => pp31(39),
		cout => pp27(40)
		);

	FA115: full_adder port map(
		a => pp18(39),
		b => pp19(39),
		cin => pp20(39),
		s => pp32(39),
		cout => pp28(40)
		);

	FA116: full_adder port map(
		a => pp8(26),
		b => pp9(24),
		cin => pp10(22),
		s => pp29(40),
		cout => pp25(41)
		);

	FA117: full_adder port map(
		a => pp11(20),
		b => pp12(18),
		cin => pp13(16),
		s => pp30(40),
		cout => pp26(41)
		);

	FA118: full_adder port map(
		a => pp14(14),
		b => pp15(12),
		cin => pp16(10),
		s => pp31(40),
		cout => pp27(41)
		);

	FA119: full_adder port map(
		a => pp17(40),
		b => pp18(40),
		cin => pp19(40),
		s => pp32(40),
		cout => pp28(41)
		);

	FA120: full_adder port map(
		a => pp7(29),
		b => pp8(27),
		cin => pp9(25),
		s => pp29(41),
		cout => pp25(42)
		);

	FA121: full_adder port map(
		a => pp10(23),
		b => pp11(21),
		cin => pp12(19),
		s => pp30(41),
		cout => pp26(42)
		);

	FA122: full_adder port map(
		a => pp13(17),
		b => pp14(15),
		cin => pp15(13),
		s => pp31(41),
		cout => pp27(42)
		);

	FA123: full_adder port map(
		a => pp16(11),
		b => pp17(41),
		cin => pp18(41),
		s => pp32(41),
		cout => pp28(42)
		);

	FA124: full_adder port map(
		a => pp6(32),
		b => pp7(30),
		cin => pp8(28),
		s => pp29(42),
		cout => pp25(43)
		);

	FA125: full_adder port map(
		a => pp9(26),
		b => pp10(24),
		cin => pp11(22),
		s => pp30(42),
		cout => pp26(43)
		);

	FA126: full_adder port map(
		a => pp12(20),
		b => pp13(18),
		cin => pp14(16),
		s => pp31(42),
		cout => pp27(43)
		);

	FA127: full_adder port map(
		a => pp15(14),
		b => pp16(12),
		cin => pp17(42),
		s => pp32(42),
		cout => pp28(43)
		);

	FA128: full_adder port map(
		a => pp5(35),
		b => pp6(33),
		cin => pp7(31),
		s => pp29(43),
		cout => pp25(44)
		);

	FA129: full_adder port map(
		a => pp8(29),
		b => pp9(27),
		cin => pp10(25),
		s => pp30(43),
		cout => pp26(44)
		);

	FA130: full_adder port map(
		a => pp11(23),
		b => pp12(21),
		cin => pp13(19),
		s => pp31(43),
		cout => pp27(44)
		);

	FA131: full_adder port map(
		a => pp14(17),
		b => pp15(15),
		cin => pp16(13),
		s => pp32(43),
		cout => pp28(44)
		);

	FA132: full_adder port map(
		a => pp5(36),
		b => pp6(34),
		cin => pp7(32),
		s => pp29(44),
		cout => pp25(45)
		);

	FA133: full_adder port map(
		a => pp8(30),
		b => pp9(28),
		cin => pp10(26),
		s => pp30(44),
		cout => pp26(45)
		);

	FA134: full_adder port map(
		a => pp11(24),
		b => pp12(22),
		cin => pp13(20),
		s => pp31(44),
		cout => pp27(45)
		);

	HA20: half_adder port map(
		a => pp14(18),
		b => pp15(16),
		s => pp32(44),
		cout => pp28(45)
		);

	FA135: full_adder port map(
		a => pp6(35),
		b => pp7(33),
		cin => pp8(31),
		s => pp29(45),
		cout => pp25(46)
		);

	FA136: full_adder port map(
		a => pp9(29),
		b => pp10(27),
		cin => pp11(25),
		s => pp30(45),
		cout => pp26(46)
		);

	FA137: full_adder port map(
		a => pp12(23),
		b => pp13(21),
		cin => pp14(19),
		s => pp31(45),
		cout => pp27(46)
		);

	FA138: full_adder port map(
		a => pp6(36),
		b => pp7(34),
		cin => pp8(32),
		s => pp28(46),
		cout => pp25(47)
		);

	FA139: full_adder port map(
		a => pp9(30),
		b => pp10(28),
		cin => pp11(26),
		s => pp29(46),
		cout => pp26(47)
		);

	HA21: half_adder port map(
		a => pp12(24),
		b => pp13(22),
		s => pp30(46),
		cout => pp27(47)
		);

	FA140: full_adder port map(
		a => pp7(35),
		b => pp8(33),
		cin => pp9(31),
		s => pp28(47),
		cout => pp25(48)
		);

	FA141: full_adder port map(
		a => pp10(29),
		b => pp11(27),
		cin => pp12(25),
		s => pp29(47),
		cout => pp26(48)
		);

	FA142: full_adder port map(
		a => pp7(36),
		b => pp8(34),
		cin => pp9(32),
		s => pp27(48),
		cout => pp25(49)
		);

	HA22: half_adder port map(
		a => pp10(30),
		b => pp11(28),
		s => pp28(48),
		cout => pp26(49)
		);

	FA143: full_adder port map(
		a => pp8(35),
		b => pp9(33),
		cin => pp10(31),
		s => pp27(49),
		cout => pp25(50)
		);

	HA23: half_adder port map(
		a => pp8(36),
		b => pp9(34),
		s => pp26(50),
		cout => pp25(51)
		);

	HA24: half_adder port map(
		a => pp0(10),
		b => pp1(10),
		s => pp33(10),
		cout => pp33(11)
		);

	HA25: half_adder port map(
		a => pp0(11),
		b => pp1(11),
		s => pp34(11),
		cout => pp33(12)
		);

	FA144: full_adder port map(
		a => pp0(12),
		b => pp1(12),
		cin => pp2(10),
		s => pp34(12),
		cout => pp33(13)
		);

	HA26: half_adder port map(
		a => pp3(8),
		b => pp4(6),
		s => pp35(12),
		cout => pp34(13)
		);

	FA145: full_adder port map(
		a => pp0(13),
		b => pp1(13),
		cin => pp2(11),
		s => pp35(13),
		cout => pp33(14)
		);

	HA27: half_adder port map(
		a => pp3(9),
		b => pp4(7),
		s => pp36(13),
		cout => pp34(14)
		);

	FA146: full_adder port map(
		a => pp0(14),
		b => pp1(14),
		cin => pp2(12),
		s => pp35(14),
		cout => pp33(15)
		);

	FA147: full_adder port map(
		a => pp3(10),
		b => pp4(8),
		cin => pp5(6),
		s => pp36(14),
		cout => pp34(15)
		);

	HA28: half_adder port map(
		a => pp6(4),
		b => pp7(2),
		s => pp37(14),
		cout => pp35(15)
		);

	FA148: full_adder port map(
		a => pp0(15),
		b => pp1(15),
		cin => pp2(13),
		s => pp36(15),
		cout => pp33(16)
		);

	FA149: full_adder port map(
		a => pp3(11),
		b => pp4(9),
		cin => pp5(7),
		s => pp37(15),
		cout => pp34(16)
		);

	HA29: half_adder port map(
		a => pp6(5),
		b => pp7(3),
		s => pp38(15),
		cout => pp35(16)
		);

	FA150: full_adder port map(
		a => pp2(14),
		b => pp3(12),
		cin => pp4(10),
		s => pp36(16),
		cout => pp33(17)
		);

	FA151: full_adder port map(
		a => pp5(8),
		b => pp6(6),
		cin => pp7(4),
		s => pp37(16),
		cout => pp34(17)
		);

	FA152: full_adder port map(
		a => pp8(2),
		b => pp9(0),
		cin => pp25(16),
		s => pp38(16),
		cout => pp35(17)
		);

	FA153: full_adder port map(
		a => pp2(15),
		b => pp3(13),
		cin => pp4(11),
		s => pp36(17),
		cout => pp33(18)
		);

	FA154: full_adder port map(
		a => pp5(9),
		b => pp6(7),
		cin => pp7(5),
		s => pp37(17),
		cout => pp34(18)
		);

	FA155: full_adder port map(
		a => pp8(3),
		b => pp25(17),
		cin => pp26(17),
		s => pp38(17),
		cout => pp35(18)
		);

	FA156: full_adder port map(
		a => pp5(10),
		b => pp6(8),
		cin => pp7(6),
		s => pp36(18),
		cout => pp33(19)
		);

	FA157: full_adder port map(
		a => pp8(4),
		b => pp9(2),
		cin => pp10(0),
		s => pp37(18),
		cout => pp34(19)
		);

	FA158: full_adder port map(
		a => pp25(18),
		b => pp26(18),
		cin => pp27(18),
		s => pp38(18),
		cout => pp35(19)
		);

	FA159: full_adder port map(
		a => pp5(11),
		b => pp6(9),
		cin => pp7(7),
		s => pp36(19),
		cout => pp33(20)
		);

	FA160: full_adder port map(
		a => pp8(5),
		b => pp9(3),
		cin => pp25(19),
		s => pp37(19),
		cout => pp34(20)
		);

	FA161: full_adder port map(
		a => pp26(19),
		b => pp27(19),
		cin => pp28(19),
		s => pp38(19),
		cout => pp35(20)
		);

	FA162: full_adder port map(
		a => pp8(6),
		b => pp9(4),
		cin => pp10(2),
		s => pp36(20),
		cout => pp33(21)
		);

	FA163: full_adder port map(
		a => pp11(0),
		b => pp25(20),
		cin => pp26(20),
		s => pp37(20),
		cout => pp34(21)
		);

	FA164: full_adder port map(
		a => pp27(20),
		b => pp28(20),
		cin => pp29(20),
		s => pp38(20),
		cout => pp35(21)
		);

	FA165: full_adder port map(
		a => pp8(7),
		b => pp9(5),
		cin => pp10(3),
		s => pp36(21),
		cout => pp33(22)
		);

	FA166: full_adder port map(
		a => pp25(21),
		b => pp26(21),
		cin => pp27(21),
		s => pp37(21),
		cout => pp34(22)
		);

	FA167: full_adder port map(
		a => pp28(21),
		b => pp29(21),
		cin => pp30(21),
		s => pp38(21),
		cout => pp35(22)
		);

	FA168: full_adder port map(
		a => pp11(2),
		b => pp12(0),
		cin => pp25(22),
		s => pp36(22),
		cout => pp33(23)
		);

	FA169: full_adder port map(
		a => pp26(22),
		b => pp27(22),
		cin => pp28(22),
		s => pp37(22),
		cout => pp34(23)
		);

	FA170: full_adder port map(
		a => pp29(22),
		b => pp30(22),
		cin => pp31(22),
		s => pp38(22),
		cout => pp35(23)
		);

	FA171: full_adder port map(
		a => pp11(3),
		b => pp25(23),
		cin => pp26(23),
		s => pp36(23),
		cout => pp33(24)
		);

	FA172: full_adder port map(
		a => pp27(23),
		b => pp28(23),
		cin => pp29(23),
		s => pp37(23),
		cout => pp34(24)
		);

	FA173: full_adder port map(
		a => pp30(23),
		b => pp31(23),
		cin => pp32(23),
		s => pp38(23),
		cout => pp35(24)
		);

	FA174: full_adder port map(
		a => pp17(24),
		b => pp25(24),
		cin => pp26(24),
		s => pp36(24),
		cout => pp33(25)
		);

	FA175: full_adder port map(
		a => pp27(24),
		b => pp28(24),
		cin => pp29(24),
		s => pp37(24),
		cout => pp34(25)
		);

	FA176: full_adder port map(
		a => pp30(24),
		b => pp31(24),
		cin => pp32(24),
		s => pp38(24),
		cout => pp35(25)
		);

	FA177: full_adder port map(
		a => pp18(25),
		b => pp25(25),
		cin => pp26(25),
		s => pp36(25),
		cout => pp33(26)
		);

	FA178: full_adder port map(
		a => pp27(25),
		b => pp28(25),
		cin => pp29(25),
		s => pp37(25),
		cout => pp34(26)
		);

	FA179: full_adder port map(
		a => pp30(25),
		b => pp31(25),
		cin => pp32(25),
		s => pp38(25),
		cout => pp35(26)
		);

	FA180: full_adder port map(
		a => pp19(26),
		b => pp25(26),
		cin => pp26(26),
		s => pp36(26),
		cout => pp33(27)
		);

	FA181: full_adder port map(
		a => pp27(26),
		b => pp28(26),
		cin => pp29(26),
		s => pp37(26),
		cout => pp34(27)
		);

	FA182: full_adder port map(
		a => pp30(26),
		b => pp31(26),
		cin => pp32(26),
		s => pp38(26),
		cout => pp35(27)
		);

	FA183: full_adder port map(
		a => pp20(27),
		b => pp25(27),
		cin => pp26(27),
		s => pp36(27),
		cout => pp33(28)
		);

	FA184: full_adder port map(
		a => pp27(27),
		b => pp28(27),
		cin => pp29(27),
		s => pp37(27),
		cout => pp34(28)
		);

	FA185: full_adder port map(
		a => pp30(27),
		b => pp31(27),
		cin => pp32(27),
		s => pp38(27),
		cout => pp35(28)
		);

	FA186: full_adder port map(
		a => pp21(28),
		b => pp25(28),
		cin => pp26(28),
		s => pp36(28),
		cout => pp33(29)
		);

	FA187: full_adder port map(
		a => pp27(28),
		b => pp28(28),
		cin => pp29(28),
		s => pp37(28),
		cout => pp34(29)
		);

	FA188: full_adder port map(
		a => pp30(28),
		b => pp31(28),
		cin => pp32(28),
		s => pp38(28),
		cout => pp35(29)
		);

	FA189: full_adder port map(
		a => pp22(29),
		b => pp25(29),
		cin => pp26(29),
		s => pp36(29),
		cout => pp33(30)
		);

	FA190: full_adder port map(
		a => pp27(29),
		b => pp28(29),
		cin => pp29(29),
		s => pp37(29),
		cout => pp34(30)
		);

	FA191: full_adder port map(
		a => pp30(29),
		b => pp31(29),
		cin => pp32(29),
		s => pp38(29),
		cout => pp35(30)
		);

	FA192: full_adder port map(
		a => pp23(30),
		b => pp25(30),
		cin => pp26(30),
		s => pp36(30),
		cout => pp33(31)
		);

	FA193: full_adder port map(
		a => pp27(30),
		b => pp28(30),
		cin => pp29(30),
		s => pp37(30),
		cout => pp34(31)
		);

	FA194: full_adder port map(
		a => pp30(30),
		b => pp31(30),
		cin => pp32(30),
		s => pp38(30),
		cout => pp35(31)
		);

	FA195: full_adder port map(
		a => pp24(31),
		b => pp25(31),
		cin => pp26(31),
		s => pp36(31),
		cout => pp33(32)
		);

	FA196: full_adder port map(
		a => pp27(31),
		b => pp28(31),
		cin => pp29(31),
		s => pp37(31),
		cout => pp34(32)
		);

	FA197: full_adder port map(
		a => pp30(31),
		b => pp31(31),
		cin => pp32(31),
		s => pp38(31),
		cout => pp35(32)
		);

	FA198: full_adder port map(
		a => pp24(32),
		b => pp25(32),
		cin => pp26(32),
		s => pp36(32),
		cout => pp33(33)
		);

	FA199: full_adder port map(
		a => pp27(32),
		b => pp28(32),
		cin => pp29(32),
		s => pp37(32),
		cout => pp34(33)
		);

	FA200: full_adder port map(
		a => pp30(32),
		b => pp31(32),
		cin => pp32(32),
		s => pp38(32),
		cout => pp35(33)
		);

	FA201: full_adder port map(
		a => pp24(33),
		b => pp25(33),
		cin => pp26(33),
		s => pp36(33),
		cout => pp33(34)
		);

	FA202: full_adder port map(
		a => pp27(33),
		b => pp28(33),
		cin => pp29(33),
		s => pp37(33),
		cout => pp34(34)
		);

	FA203: full_adder port map(
		a => pp30(33),
		b => pp31(33),
		cin => pp32(33),
		s => pp38(33),
		cout => pp35(34)
		);

	FA204: full_adder port map(
		a => pp24(34),
		b => pp25(34),
		cin => pp26(34),
		s => pp36(34),
		cout => pp33(35)
		);

	FA205: full_adder port map(
		a => pp27(34),
		b => pp28(34),
		cin => pp29(34),
		s => pp37(34),
		cout => pp34(35)
		);

	FA206: full_adder port map(
		a => pp30(34),
		b => pp31(34),
		cin => pp32(34),
		s => pp38(34),
		cout => pp35(35)
		);

	FA207: full_adder port map(
		a => pp24(35),
		b => pp25(35),
		cin => pp26(35),
		s => pp36(35),
		cout => pp33(36)
		);

	FA208: full_adder port map(
		a => pp27(35),
		b => pp28(35),
		cin => pp29(35),
		s => pp37(35),
		cout => pp34(36)
		);

	FA209: full_adder port map(
		a => pp30(35),
		b => pp31(35),
		cin => pp32(35),
		s => pp38(35),
		cout => pp35(36)
		);

	FA210: full_adder port map(
		a => pp24(36),
		b => pp25(36),
		cin => pp26(36),
		s => pp36(36),
		cout => pp33(37)
		);

	FA211: full_adder port map(
		a => pp27(36),
		b => pp28(36),
		cin => pp29(36),
		s => pp37(36),
		cout => pp34(37)
		);

	FA212: full_adder port map(
		a => pp30(36),
		b => pp31(36),
		cin => pp32(36),
		s => pp38(36),
		cout => pp35(37)
		);

	FA213: full_adder port map(
		a => pp23(37),
		b => pp25(37),
		cin => pp26(37),
		s => pp36(37),
		cout => pp33(38)
		);

	FA214: full_adder port map(
		a => pp27(37),
		b => pp28(37),
		cin => pp29(37),
		s => pp37(37),
		cout => pp34(38)
		);

	FA215: full_adder port map(
		a => pp30(37),
		b => pp31(37),
		cin => pp32(37),
		s => pp38(37),
		cout => pp35(38)
		);

	FA216: full_adder port map(
		a => pp22(38),
		b => pp25(38),
		cin => pp26(38),
		s => pp36(38),
		cout => pp33(39)
		);

	FA217: full_adder port map(
		a => pp27(38),
		b => pp28(38),
		cin => pp29(38),
		s => pp37(38),
		cout => pp34(39)
		);

	FA218: full_adder port map(
		a => pp30(38),
		b => pp31(38),
		cin => pp32(38),
		s => pp38(38),
		cout => pp35(39)
		);

	FA219: full_adder port map(
		a => pp21(39),
		b => pp25(39),
		cin => pp26(39),
		s => pp36(39),
		cout => pp33(40)
		);

	FA220: full_adder port map(
		a => pp27(39),
		b => pp28(39),
		cin => pp29(39),
		s => pp37(39),
		cout => pp34(40)
		);

	FA221: full_adder port map(
		a => pp30(39),
		b => pp31(39),
		cin => pp32(39),
		s => pp38(39),
		cout => pp35(40)
		);

	FA222: full_adder port map(
		a => pp20(40),
		b => pp25(40),
		cin => pp26(40),
		s => pp36(40),
		cout => pp33(41)
		);

	FA223: full_adder port map(
		a => pp27(40),
		b => pp28(40),
		cin => pp29(40),
		s => pp37(40),
		cout => pp34(41)
		);

	FA224: full_adder port map(
		a => pp30(40),
		b => pp31(40),
		cin => pp32(40),
		s => pp38(40),
		cout => pp35(41)
		);

	FA225: full_adder port map(
		a => pp19(41),
		b => pp25(41),
		cin => pp26(41),
		s => pp36(41),
		cout => pp33(42)
		);

	FA226: full_adder port map(
		a => pp27(41),
		b => pp28(41),
		cin => pp29(41),
		s => pp37(41),
		cout => pp34(42)
		);

	FA227: full_adder port map(
		a => pp30(41),
		b => pp31(41),
		cin => pp32(41),
		s => pp38(41),
		cout => pp35(42)
		);

	FA228: full_adder port map(
		a => pp18(42),
		b => pp25(42),
		cin => pp26(42),
		s => pp36(42),
		cout => pp33(43)
		);

	FA229: full_adder port map(
		a => pp27(42),
		b => pp28(42),
		cin => pp29(42),
		s => pp37(42),
		cout => pp34(43)
		);

	FA230: full_adder port map(
		a => pp30(42),
		b => pp31(42),
		cin => pp32(42),
		s => pp38(42),
		cout => pp35(43)
		);

	FA231: full_adder port map(
		a => pp17(43),
		b => pp25(43),
		cin => pp26(43),
		s => pp36(43),
		cout => pp33(44)
		);

	FA232: full_adder port map(
		a => pp27(43),
		b => pp28(43),
		cin => pp29(43),
		s => pp37(43),
		cout => pp34(44)
		);

	FA233: full_adder port map(
		a => pp30(43),
		b => pp31(43),
		cin => pp32(43),
		s => pp38(43),
		cout => pp35(44)
		);

	FA234: full_adder port map(
		a => pp16(14),
		b => pp25(44),
		cin => pp26(44),
		s => pp36(44),
		cout => pp33(45)
		);

	FA235: full_adder port map(
		a => pp27(44),
		b => pp28(44),
		cin => pp29(44),
		s => pp37(44),
		cout => pp34(45)
		);

	FA236: full_adder port map(
		a => pp30(44),
		b => pp31(44),
		cin => pp32(44),
		s => pp38(44),
		cout => pp35(45)
		);

	FA237: full_adder port map(
		a => pp15(17),
		b => pp16(15),
		cin => pp25(45),
		s => pp36(45),
		cout => pp33(46)
		);

	FA238: full_adder port map(
		a => pp26(45),
		b => pp27(45),
		cin => pp28(45),
		s => pp37(45),
		cout => pp34(46)
		);

	FA239: full_adder port map(
		a => pp29(45),
		b => pp30(45),
		cin => pp31(45),
		s => pp38(45),
		cout => pp35(46)
		);

	FA240: full_adder port map(
		a => pp14(20),
		b => pp15(18),
		cin => pp16(16),
		s => pp36(46),
		cout => pp33(47)
		);

	FA241: full_adder port map(
		a => pp25(46),
		b => pp26(46),
		cin => pp27(46),
		s => pp37(46),
		cout => pp34(47)
		);

	FA242: full_adder port map(
		a => pp28(46),
		b => pp29(46),
		cin => pp30(46),
		s => pp38(46),
		cout => pp35(47)
		);

	FA243: full_adder port map(
		a => pp13(23),
		b => pp14(21),
		cin => pp15(19),
		s => pp36(47),
		cout => pp33(48)
		);

	FA244: full_adder port map(
		a => pp16(17),
		b => pp25(47),
		cin => pp26(47),
		s => pp37(47),
		cout => pp34(48)
		);

	FA245: full_adder port map(
		a => pp27(47),
		b => pp28(47),
		cin => pp29(47),
		s => pp38(47),
		cout => pp35(48)
		);

	FA246: full_adder port map(
		a => pp12(26),
		b => pp13(24),
		cin => pp14(22),
		s => pp36(48),
		cout => pp33(49)
		);

	FA247: full_adder port map(
		a => pp15(20),
		b => pp16(18),
		cin => pp25(48),
		s => pp37(48),
		cout => pp34(49)
		);

	FA248: full_adder port map(
		a => pp26(48),
		b => pp27(48),
		cin => pp28(48),
		s => pp38(48),
		cout => pp35(49)
		);

	FA249: full_adder port map(
		a => pp11(29),
		b => pp12(27),
		cin => pp13(25),
		s => pp36(49),
		cout => pp33(50)
		);

	FA250: full_adder port map(
		a => pp14(23),
		b => pp15(21),
		cin => pp16(19),
		s => pp37(49),
		cout => pp34(50)
		);

	FA251: full_adder port map(
		a => pp25(49),
		b => pp26(49),
		cin => pp27(49),
		s => pp38(49),
		cout => pp35(50)
		);

	FA252: full_adder port map(
		a => pp10(32),
		b => pp11(30),
		cin => pp12(28),
		s => pp36(50),
		cout => pp33(51)
		);

	FA253: full_adder port map(
		a => pp13(26),
		b => pp14(24),
		cin => pp15(22),
		s => pp37(50),
		cout => pp34(51)
		);

	FA254: full_adder port map(
		a => pp16(20),
		b => pp25(50),
		cin => pp26(50),
		s => pp38(50),
		cout => pp35(51)
		);

	FA255: full_adder port map(
		a => pp9(35),
		b => pp10(33),
		cin => pp11(31),
		s => pp36(51),
		cout => pp33(52)
		);

	FA256: full_adder port map(
		a => pp12(29),
		b => pp13(27),
		cin => pp14(25),
		s => pp37(51),
		cout => pp34(52)
		);

	FA257: full_adder port map(
		a => pp15(23),
		b => pp16(21),
		cin => pp25(51),
		s => pp38(51),
		cout => pp35(52)
		);

	FA258: full_adder port map(
		a => pp9(36),
		b => pp10(34),
		cin => pp11(32),
		s => pp36(52),
		cout => pp33(53)
		);

	FA259: full_adder port map(
		a => pp12(30),
		b => pp13(28),
		cin => pp14(26),
		s => pp37(52),
		cout => pp34(53)
		);

	HA30: half_adder port map(
		a => pp15(24),
		b => pp16(22),
		s => pp38(52),
		cout => pp35(53)
		);

	FA260: full_adder port map(
		a => pp10(35),
		b => pp11(33),
		cin => pp12(31),
		s => pp36(53),
		cout => pp33(54)
		);

	FA261: full_adder port map(
		a => pp13(29),
		b => pp14(27),
		cin => pp15(25),
		s => pp37(53),
		cout => pp34(54)
		);

	FA262: full_adder port map(
		a => pp10(36),
		b => pp11(34),
		cin => pp12(32),
		s => pp35(54),
		cout => pp33(55)
		);

	HA31: half_adder port map(
		a => pp13(30),
		b => pp14(28),
		s => pp36(54),
		cout => pp34(55)
		);

	FA263: full_adder port map(
		a => pp11(35),
		b => pp12(33),
		cin => pp13(31),
		s => pp35(55),
		cout => pp33(56)
		);

	HA32: half_adder port map(
		a => pp11(36),
		b => pp12(34),
		s => pp34(56),
		cout => pp33(57)
		);

	HA33: half_adder port map(
		a => pp0(6),
		b => pp1(6),
		s => pp39(6),
		cout => pp39(7)
		);

	HA34: half_adder port map(
		a => pp0(7),
		b => pp1(7),
		s => pp40(7),
		cout => pp39(8)
		);

	FA264: full_adder port map(
		a => pp0(8),
		b => pp1(8),
		cin => pp2(6),
		s => pp40(8),
		cout => pp39(9)
		);

	HA35: half_adder port map(
		a => pp3(4),
		b => pp4(2),
		s => pp41(8),
		cout => pp40(9)
		);

	FA265: full_adder port map(
		a => pp0(9),
		b => pp1(9),
		cin => pp2(7),
		s => pp41(9),
		cout => pp39(10)
		);

	HA36: half_adder port map(
		a => pp3(5),
		b => pp4(3),
		s => pp42(9),
		cout => pp40(10)
		);

	FA266: full_adder port map(
		a => pp2(8),
		b => pp3(6),
		cin => pp4(4),
		s => pp41(10),
		cout => pp39(11)
		);

	FA267: full_adder port map(
		a => pp5(2),
		b => pp6(0),
		cin => pp33(10),
		s => pp42(10),
		cout => pp40(11)
		);

	FA268: full_adder port map(
		a => pp2(9),
		b => pp3(7),
		cin => pp4(5),
		s => pp41(11),
		cout => pp39(12)
		);

	FA269: full_adder port map(
		a => pp5(3),
		b => pp33(11),
		cin => pp34(11),
		s => pp42(11),
		cout => pp40(12)
		);

	FA270: full_adder port map(
		a => pp5(4),
		b => pp6(2),
		cin => pp7(0),
		s => pp41(12),
		cout => pp39(13)
		);

	FA271: full_adder port map(
		a => pp33(12),
		b => pp34(12),
		cin => pp35(12),
		s => pp42(12),
		cout => pp40(13)
		);

	FA272: full_adder port map(
		a => pp5(5),
		b => pp6(3),
		cin => pp33(13),
		s => pp41(13),
		cout => pp39(14)
		);

	FA273: full_adder port map(
		a => pp34(13),
		b => pp35(13),
		cin => pp36(13),
		s => pp42(13),
		cout => pp40(14)
		);

	FA274: full_adder port map(
		a => pp8(0),
		b => pp33(14),
		cin => pp34(14),
		s => pp41(14),
		cout => pp39(15)
		);

	FA275: full_adder port map(
		a => pp35(14),
		b => pp36(14),
		cin => pp37(14),
		s => pp42(14),
		cout => pp40(15)
		);

	FA276: full_adder port map(
		a => pp33(15),
		b => pp34(15),
		cin => pp35(15),
		s => pp41(15),
		cout => pp39(16)
		);

	FA277: full_adder port map(
		a => pp36(15),
		b => pp37(15),
		cin => pp38(15),
		s => pp42(15),
		cout => pp40(16)
		);

	FA278: full_adder port map(
		a => pp33(16),
		b => pp34(16),
		cin => pp35(16),
		s => pp41(16),
		cout => pp39(17)
		);

	FA279: full_adder port map(
		a => pp36(16),
		b => pp37(16),
		cin => pp38(16),
		s => pp42(16),
		cout => pp40(17)
		);

	FA280: full_adder port map(
		a => pp33(17),
		b => pp34(17),
		cin => pp35(17),
		s => pp41(17),
		cout => pp39(18)
		);

	FA281: full_adder port map(
		a => pp36(17),
		b => pp37(17),
		cin => pp38(17),
		s => pp42(17),
		cout => pp40(18)
		);

	FA282: full_adder port map(
		a => pp33(18),
		b => pp34(18),
		cin => pp35(18),
		s => pp41(18),
		cout => pp39(19)
		);

	FA283: full_adder port map(
		a => pp36(18),
		b => pp37(18),
		cin => pp38(18),
		s => pp42(18),
		cout => pp40(19)
		);

	FA284: full_adder port map(
		a => pp33(19),
		b => pp34(19),
		cin => pp35(19),
		s => pp41(19),
		cout => pp39(20)
		);

	FA285: full_adder port map(
		a => pp36(19),
		b => pp37(19),
		cin => pp38(19),
		s => pp42(19),
		cout => pp40(20)
		);

	FA286: full_adder port map(
		a => pp33(20),
		b => pp34(20),
		cin => pp35(20),
		s => pp41(20),
		cout => pp39(21)
		);

	FA287: full_adder port map(
		a => pp36(20),
		b => pp37(20),
		cin => pp38(20),
		s => pp42(20),
		cout => pp40(21)
		);

	FA288: full_adder port map(
		a => pp33(21),
		b => pp34(21),
		cin => pp35(21),
		s => pp41(21),
		cout => pp39(22)
		);

	FA289: full_adder port map(
		a => pp36(21),
		b => pp37(21),
		cin => pp38(21),
		s => pp42(21),
		cout => pp40(22)
		);

	FA290: full_adder port map(
		a => pp33(22),
		b => pp34(22),
		cin => pp35(22),
		s => pp41(22),
		cout => pp39(23)
		);

	FA291: full_adder port map(
		a => pp36(22),
		b => pp37(22),
		cin => pp38(22),
		s => pp42(22),
		cout => pp40(23)
		);

	FA292: full_adder port map(
		a => pp33(23),
		b => pp34(23),
		cin => pp35(23),
		s => pp41(23),
		cout => pp39(24)
		);

	FA293: full_adder port map(
		a => pp36(23),
		b => pp37(23),
		cin => pp38(23),
		s => pp42(23),
		cout => pp40(24)
		);

	FA294: full_adder port map(
		a => pp33(24),
		b => pp34(24),
		cin => pp35(24),
		s => pp41(24),
		cout => pp39(25)
		);

	FA295: full_adder port map(
		a => pp36(24),
		b => pp37(24),
		cin => pp38(24),
		s => pp42(24),
		cout => pp40(25)
		);

	FA296: full_adder port map(
		a => pp33(25),
		b => pp34(25),
		cin => pp35(25),
		s => pp41(25),
		cout => pp39(26)
		);

	FA297: full_adder port map(
		a => pp36(25),
		b => pp37(25),
		cin => pp38(25),
		s => pp42(25),
		cout => pp40(26)
		);

	FA298: full_adder port map(
		a => pp33(26),
		b => pp34(26),
		cin => pp35(26),
		s => pp41(26),
		cout => pp39(27)
		);

	FA299: full_adder port map(
		a => pp36(26),
		b => pp37(26),
		cin => pp38(26),
		s => pp42(26),
		cout => pp40(27)
		);

	FA300: full_adder port map(
		a => pp33(27),
		b => pp34(27),
		cin => pp35(27),
		s => pp41(27),
		cout => pp39(28)
		);

	FA301: full_adder port map(
		a => pp36(27),
		b => pp37(27),
		cin => pp38(27),
		s => pp42(27),
		cout => pp40(28)
		);

	FA302: full_adder port map(
		a => pp33(28),
		b => pp34(28),
		cin => pp35(28),
		s => pp41(28),
		cout => pp39(29)
		);

	FA303: full_adder port map(
		a => pp36(28),
		b => pp37(28),
		cin => pp38(28),
		s => pp42(28),
		cout => pp40(29)
		);

	FA304: full_adder port map(
		a => pp33(29),
		b => pp34(29),
		cin => pp35(29),
		s => pp41(29),
		cout => pp39(30)
		);

	FA305: full_adder port map(
		a => pp36(29),
		b => pp37(29),
		cin => pp38(29),
		s => pp42(29),
		cout => pp40(30)
		);

	FA306: full_adder port map(
		a => pp33(30),
		b => pp34(30),
		cin => pp35(30),
		s => pp41(30),
		cout => pp39(31)
		);

	FA307: full_adder port map(
		a => pp36(30),
		b => pp37(30),
		cin => pp38(30),
		s => pp42(30),
		cout => pp40(31)
		);

	FA308: full_adder port map(
		a => pp33(31),
		b => pp34(31),
		cin => pp35(31),
		s => pp41(31),
		cout => pp39(32)
		);

	FA309: full_adder port map(
		a => pp36(31),
		b => pp37(31),
		cin => pp38(31),
		s => pp42(31),
		cout => pp40(32)
		);

	FA310: full_adder port map(
		a => pp33(32),
		b => pp34(32),
		cin => pp35(32),
		s => pp41(32),
		cout => pp39(33)
		);

	FA311: full_adder port map(
		a => pp36(32),
		b => pp37(32),
		cin => pp38(32),
		s => pp42(32),
		cout => pp40(33)
		);

	FA312: full_adder port map(
		a => pp33(33),
		b => pp34(33),
		cin => pp35(33),
		s => pp41(33),
		cout => pp39(34)
		);

	FA313: full_adder port map(
		a => pp36(33),
		b => pp37(33),
		cin => pp38(33),
		s => pp42(33),
		cout => pp40(34)
		);

	FA314: full_adder port map(
		a => pp33(34),
		b => pp34(34),
		cin => pp35(34),
		s => pp41(34),
		cout => pp39(35)
		);

	FA315: full_adder port map(
		a => pp36(34),
		b => pp37(34),
		cin => pp38(34),
		s => pp42(34),
		cout => pp40(35)
		);

	FA316: full_adder port map(
		a => pp33(35),
		b => pp34(35),
		cin => pp35(35),
		s => pp41(35),
		cout => pp39(36)
		);

	FA317: full_adder port map(
		a => pp36(35),
		b => pp37(35),
		cin => pp38(35),
		s => pp42(35),
		cout => pp40(36)
		);

	FA318: full_adder port map(
		a => pp33(36),
		b => pp34(36),
		cin => pp35(36),
		s => pp41(36),
		cout => pp39(37)
		);

	FA319: full_adder port map(
		a => pp36(36),
		b => pp37(36),
		cin => pp38(36),
		s => pp42(36),
		cout => pp40(37)
		);

	FA320: full_adder port map(
		a => pp33(37),
		b => pp34(37),
		cin => pp35(37),
		s => pp41(37),
		cout => pp39(38)
		);

	FA321: full_adder port map(
		a => pp36(37),
		b => pp37(37),
		cin => pp38(37),
		s => pp42(37),
		cout => pp40(38)
		);

	FA322: full_adder port map(
		a => pp33(38),
		b => pp34(38),
		cin => pp35(38),
		s => pp41(38),
		cout => pp39(39)
		);

	FA323: full_adder port map(
		a => pp36(38),
		b => pp37(38),
		cin => pp38(38),
		s => pp42(38),
		cout => pp40(39)
		);

	FA324: full_adder port map(
		a => pp33(39),
		b => pp34(39),
		cin => pp35(39),
		s => pp41(39),
		cout => pp39(40)
		);

	FA325: full_adder port map(
		a => pp36(39),
		b => pp37(39),
		cin => pp38(39),
		s => pp42(39),
		cout => pp40(40)
		);

	FA326: full_adder port map(
		a => pp33(40),
		b => pp34(40),
		cin => pp35(40),
		s => pp41(40),
		cout => pp39(41)
		);

	FA327: full_adder port map(
		a => pp36(40),
		b => pp37(40),
		cin => pp38(40),
		s => pp42(40),
		cout => pp40(41)
		);

	FA328: full_adder port map(
		a => pp33(41),
		b => pp34(41),
		cin => pp35(41),
		s => pp41(41),
		cout => pp39(42)
		);

	FA329: full_adder port map(
		a => pp36(41),
		b => pp37(41),
		cin => pp38(41),
		s => pp42(41),
		cout => pp40(42)
		);

	FA330: full_adder port map(
		a => pp33(42),
		b => pp34(42),
		cin => pp35(42),
		s => pp41(42),
		cout => pp39(43)
		);

	FA331: full_adder port map(
		a => pp36(42),
		b => pp37(42),
		cin => pp38(42),
		s => pp42(42),
		cout => pp40(43)
		);

	FA332: full_adder port map(
		a => pp33(43),
		b => pp34(43),
		cin => pp35(43),
		s => pp41(43),
		cout => pp39(44)
		);

	FA333: full_adder port map(
		a => pp36(43),
		b => pp37(43),
		cin => pp38(43),
		s => pp42(43),
		cout => pp40(44)
		);

	FA334: full_adder port map(
		a => pp33(44),
		b => pp34(44),
		cin => pp35(44),
		s => pp41(44),
		cout => pp39(45)
		);

	FA335: full_adder port map(
		a => pp36(44),
		b => pp37(44),
		cin => pp38(44),
		s => pp42(44),
		cout => pp40(45)
		);

	FA336: full_adder port map(
		a => pp33(45),
		b => pp34(45),
		cin => pp35(45),
		s => pp41(45),
		cout => pp39(46)
		);

	FA337: full_adder port map(
		a => pp36(45),
		b => pp37(45),
		cin => pp38(45),
		s => pp42(45),
		cout => pp40(46)
		);

	FA338: full_adder port map(
		a => pp33(46),
		b => pp34(46),
		cin => pp35(46),
		s => pp41(46),
		cout => pp39(47)
		);

	FA339: full_adder port map(
		a => pp36(46),
		b => pp37(46),
		cin => pp38(46),
		s => pp42(46),
		cout => pp40(47)
		);

	FA340: full_adder port map(
		a => pp33(47),
		b => pp34(47),
		cin => pp35(47),
		s => pp41(47),
		cout => pp39(48)
		);

	FA341: full_adder port map(
		a => pp36(47),
		b => pp37(47),
		cin => pp38(47),
		s => pp42(47),
		cout => pp40(48)
		);

	FA342: full_adder port map(
		a => pp33(48),
		b => pp34(48),
		cin => pp35(48),
		s => pp41(48),
		cout => pp39(49)
		);

	FA343: full_adder port map(
		a => pp36(48),
		b => pp37(48),
		cin => pp38(48),
		s => pp42(48),
		cout => pp40(49)
		);

	FA344: full_adder port map(
		a => pp33(49),
		b => pp34(49),
		cin => pp35(49),
		s => pp41(49),
		cout => pp39(50)
		);

	FA345: full_adder port map(
		a => pp36(49),
		b => pp37(49),
		cin => pp38(49),
		s => pp42(49),
		cout => pp40(50)
		);

	FA346: full_adder port map(
		a => pp33(50),
		b => pp34(50),
		cin => pp35(50),
		s => pp41(50),
		cout => pp39(51)
		);

	FA347: full_adder port map(
		a => pp36(50),
		b => pp37(50),
		cin => pp38(50),
		s => pp42(50),
		cout => pp40(51)
		);

	FA348: full_adder port map(
		a => pp33(51),
		b => pp34(51),
		cin => pp35(51),
		s => pp41(51),
		cout => pp39(52)
		);

	FA349: full_adder port map(
		a => pp36(51),
		b => pp37(51),
		cin => pp38(51),
		s => pp42(51),
		cout => pp40(52)
		);

	FA350: full_adder port map(
		a => pp33(52),
		b => pp34(52),
		cin => pp35(52),
		s => pp41(52),
		cout => pp39(53)
		);

	FA351: full_adder port map(
		a => pp36(52),
		b => pp37(52),
		cin => pp38(52),
		s => pp42(52),
		cout => pp40(53)
		);

	FA352: full_adder port map(
		a => pp16(23),
		b => pp33(53),
		cin => pp34(53),
		s => pp41(53),
		cout => pp39(54)
		);

	FA353: full_adder port map(
		a => pp35(53),
		b => pp36(53),
		cin => pp37(53),
		s => pp42(53),
		cout => pp40(54)
		);

	FA354: full_adder port map(
		a => pp15(26),
		b => pp16(24),
		cin => pp33(54),
		s => pp41(54),
		cout => pp39(55)
		);

	FA355: full_adder port map(
		a => pp34(54),
		b => pp35(54),
		cin => pp36(54),
		s => pp42(54),
		cout => pp40(55)
		);

	FA356: full_adder port map(
		a => pp14(29),
		b => pp15(27),
		cin => pp16(25),
		s => pp41(55),
		cout => pp39(56)
		);

	FA357: full_adder port map(
		a => pp33(55),
		b => pp34(55),
		cin => pp35(55),
		s => pp42(55),
		cout => pp40(56)
		);

	FA358: full_adder port map(
		a => pp13(32),
		b => pp14(30),
		cin => pp15(28),
		s => pp41(56),
		cout => pp39(57)
		);

	FA359: full_adder port map(
		a => pp16(26),
		b => pp33(56),
		cin => pp34(56),
		s => pp42(56),
		cout => pp40(57)
		);

	FA360: full_adder port map(
		a => pp12(35),
		b => pp13(33),
		cin => pp14(31),
		s => pp41(57),
		cout => pp39(58)
		);

	FA361: full_adder port map(
		a => pp15(29),
		b => pp16(27),
		cin => pp33(57),
		s => pp42(57),
		cout => pp40(58)
		);

	FA362: full_adder port map(
		a => pp12(36),
		b => pp13(34),
		cin => pp14(32),
		s => pp41(58),
		cout => pp39(59)
		);

	HA37: half_adder port map(
		a => pp15(30),
		b => pp16(28),
		s => pp42(58),
		cout => pp40(59)
		);

	FA363: full_adder port map(
		a => pp13(35),
		b => pp14(33),
		cin => pp15(31),
		s => pp41(59),
		cout => pp39(60)
		);

	HA38: half_adder port map(
		a => pp13(36),
		b => pp14(34),
		s => pp40(60),
		cout => pp39(61)
		);

	HA39: half_adder port map(
		a => pp0(4),
		b => pp1(4),
		s => pp43(4),
		cout => pp43(5)
		);

	HA40: half_adder port map(
		a => pp0(5),
		b => pp1(5),
		s => pp44(5),
		cout => pp43(6)
		);

	FA364: full_adder port map(
		a => pp2(4),
		b => pp3(2),
		cin => pp4(0),
		s => pp44(6),
		cout => pp43(7)
		);

	FA365: full_adder port map(
		a => pp2(5),
		b => pp3(3),
		cin => pp39(7),
		s => pp44(7),
		cout => pp43(8)
		);

	FA366: full_adder port map(
		a => pp5(0),
		b => pp39(8),
		cin => pp40(8),
		s => pp44(8),
		cout => pp43(9)
		);

	FA367: full_adder port map(
		a => pp39(9),
		b => pp40(9),
		cin => pp41(9),
		s => pp44(9),
		cout => pp43(10)
		);

	FA368: full_adder port map(
		a => pp39(10),
		b => pp40(10),
		cin => pp41(10),
		s => pp44(10),
		cout => pp43(11)
		);

	FA369: full_adder port map(
		a => pp39(11),
		b => pp40(11),
		cin => pp41(11),
		s => pp44(11),
		cout => pp43(12)
		);

	FA370: full_adder port map(
		a => pp39(12),
		b => pp40(12),
		cin => pp41(12),
		s => pp44(12),
		cout => pp43(13)
		);

	FA371: full_adder port map(
		a => pp39(13),
		b => pp40(13),
		cin => pp41(13),
		s => pp44(13),
		cout => pp43(14)
		);

	FA372: full_adder port map(
		a => pp39(14),
		b => pp40(14),
		cin => pp41(14),
		s => pp44(14),
		cout => pp43(15)
		);

	FA373: full_adder port map(
		a => pp39(15),
		b => pp40(15),
		cin => pp41(15),
		s => pp44(15),
		cout => pp43(16)
		);

	FA374: full_adder port map(
		a => pp39(16),
		b => pp40(16),
		cin => pp41(16),
		s => pp44(16),
		cout => pp43(17)
		);

	FA375: full_adder port map(
		a => pp39(17),
		b => pp40(17),
		cin => pp41(17),
		s => pp44(17),
		cout => pp43(18)
		);

	FA376: full_adder port map(
		a => pp39(18),
		b => pp40(18),
		cin => pp41(18),
		s => pp44(18),
		cout => pp43(19)
		);

	FA377: full_adder port map(
		a => pp39(19),
		b => pp40(19),
		cin => pp41(19),
		s => pp44(19),
		cout => pp43(20)
		);

	FA378: full_adder port map(
		a => pp39(20),
		b => pp40(20),
		cin => pp41(20),
		s => pp44(20),
		cout => pp43(21)
		);

	FA379: full_adder port map(
		a => pp39(21),
		b => pp40(21),
		cin => pp41(21),
		s => pp44(21),
		cout => pp43(22)
		);

	FA380: full_adder port map(
		a => pp39(22),
		b => pp40(22),
		cin => pp41(22),
		s => pp44(22),
		cout => pp43(23)
		);

	FA381: full_adder port map(
		a => pp39(23),
		b => pp40(23),
		cin => pp41(23),
		s => pp44(23),
		cout => pp43(24)
		);

	FA382: full_adder port map(
		a => pp39(24),
		b => pp40(24),
		cin => pp41(24),
		s => pp44(24),
		cout => pp43(25)
		);

	FA383: full_adder port map(
		a => pp39(25),
		b => pp40(25),
		cin => pp41(25),
		s => pp44(25),
		cout => pp43(26)
		);

	FA384: full_adder port map(
		a => pp39(26),
		b => pp40(26),
		cin => pp41(26),
		s => pp44(26),
		cout => pp43(27)
		);

	FA385: full_adder port map(
		a => pp39(27),
		b => pp40(27),
		cin => pp41(27),
		s => pp44(27),
		cout => pp43(28)
		);

	FA386: full_adder port map(
		a => pp39(28),
		b => pp40(28),
		cin => pp41(28),
		s => pp44(28),
		cout => pp43(29)
		);

	FA387: full_adder port map(
		a => pp39(29),
		b => pp40(29),
		cin => pp41(29),
		s => pp44(29),
		cout => pp43(30)
		);

	FA388: full_adder port map(
		a => pp39(30),
		b => pp40(30),
		cin => pp41(30),
		s => pp44(30),
		cout => pp43(31)
		);

	FA389: full_adder port map(
		a => pp39(31),
		b => pp40(31),
		cin => pp41(31),
		s => pp44(31),
		cout => pp43(32)
		);

	FA390: full_adder port map(
		a => pp39(32),
		b => pp40(32),
		cin => pp41(32),
		s => pp44(32),
		cout => pp43(33)
		);

	FA391: full_adder port map(
		a => pp39(33),
		b => pp40(33),
		cin => pp41(33),
		s => pp44(33),
		cout => pp43(34)
		);

	FA392: full_adder port map(
		a => pp39(34),
		b => pp40(34),
		cin => pp41(34),
		s => pp44(34),
		cout => pp43(35)
		);

	FA393: full_adder port map(
		a => pp39(35),
		b => pp40(35),
		cin => pp41(35),
		s => pp44(35),
		cout => pp43(36)
		);

	FA394: full_adder port map(
		a => pp39(36),
		b => pp40(36),
		cin => pp41(36),
		s => pp44(36),
		cout => pp43(37)
		);

	FA395: full_adder port map(
		a => pp39(37),
		b => pp40(37),
		cin => pp41(37),
		s => pp44(37),
		cout => pp43(38)
		);

	FA396: full_adder port map(
		a => pp39(38),
		b => pp40(38),
		cin => pp41(38),
		s => pp44(38),
		cout => pp43(39)
		);

	FA397: full_adder port map(
		a => pp39(39),
		b => pp40(39),
		cin => pp41(39),
		s => pp44(39),
		cout => pp43(40)
		);

	FA398: full_adder port map(
		a => pp39(40),
		b => pp40(40),
		cin => pp41(40),
		s => pp44(40),
		cout => pp43(41)
		);

	FA399: full_adder port map(
		a => pp39(41),
		b => pp40(41),
		cin => pp41(41),
		s => pp44(41),
		cout => pp43(42)
		);

	FA400: full_adder port map(
		a => pp39(42),
		b => pp40(42),
		cin => pp41(42),
		s => pp44(42),
		cout => pp43(43)
		);

	FA401: full_adder port map(
		a => pp39(43),
		b => pp40(43),
		cin => pp41(43),
		s => pp44(43),
		cout => pp43(44)
		);

	FA402: full_adder port map(
		a => pp39(44),
		b => pp40(44),
		cin => pp41(44),
		s => pp44(44),
		cout => pp43(45)
		);

	FA403: full_adder port map(
		a => pp39(45),
		b => pp40(45),
		cin => pp41(45),
		s => pp44(45),
		cout => pp43(46)
		);

	FA404: full_adder port map(
		a => pp39(46),
		b => pp40(46),
		cin => pp41(46),
		s => pp44(46),
		cout => pp43(47)
		);

	FA405: full_adder port map(
		a => pp39(47),
		b => pp40(47),
		cin => pp41(47),
		s => pp44(47),
		cout => pp43(48)
		);

	FA406: full_adder port map(
		a => pp39(48),
		b => pp40(48),
		cin => pp41(48),
		s => pp44(48),
		cout => pp43(49)
		);

	FA407: full_adder port map(
		a => pp39(49),
		b => pp40(49),
		cin => pp41(49),
		s => pp44(49),
		cout => pp43(50)
		);

	FA408: full_adder port map(
		a => pp39(50),
		b => pp40(50),
		cin => pp41(50),
		s => pp44(50),
		cout => pp43(51)
		);

	FA409: full_adder port map(
		a => pp39(51),
		b => pp40(51),
		cin => pp41(51),
		s => pp44(51),
		cout => pp43(52)
		);

	FA410: full_adder port map(
		a => pp39(52),
		b => pp40(52),
		cin => pp41(52),
		s => pp44(52),
		cout => pp43(53)
		);

	FA411: full_adder port map(
		a => pp39(53),
		b => pp40(53),
		cin => pp41(53),
		s => pp44(53),
		cout => pp43(54)
		);

	FA412: full_adder port map(
		a => pp39(54),
		b => pp40(54),
		cin => pp41(54),
		s => pp44(54),
		cout => pp43(55)
		);

	FA413: full_adder port map(
		a => pp39(55),
		b => pp40(55),
		cin => pp41(55),
		s => pp44(55),
		cout => pp43(56)
		);

	FA414: full_adder port map(
		a => pp39(56),
		b => pp40(56),
		cin => pp41(56),
		s => pp44(56),
		cout => pp43(57)
		);

	FA415: full_adder port map(
		a => pp39(57),
		b => pp40(57),
		cin => pp41(57),
		s => pp44(57),
		cout => pp43(58)
		);

	FA416: full_adder port map(
		a => pp39(58),
		b => pp40(58),
		cin => pp41(58),
		s => pp44(58),
		cout => pp43(59)
		);

	FA417: full_adder port map(
		a => pp16(29),
		b => pp39(59),
		cin => pp40(59),
		s => pp44(59),
		cout => pp43(60)
		);

	FA418: full_adder port map(
		a => pp15(32),
		b => pp16(30),
		cin => pp39(60),
		s => pp44(60),
		cout => pp43(61)
		);

	FA419: full_adder port map(
		a => pp14(35),
		b => pp15(33),
		cin => pp16(31),
		s => pp44(61),
		cout => pp43(62)
		);

	HA41: half_adder port map(
		a => pp14(36),
		b => pp15(34),
		s => pp44(62),
		cout => pp43(63)
		);

	HA42: half_adder port map(
		a => pp0(2),
		b => pp1(2),
		s => pp45(2),
		cout => pp45(3)
		);

	HA43: half_adder port map(
		a => pp0(3),
		b => pp1(3),
		s => pp46(3),
		cout => pp45(4)
		);

	FA420: full_adder port map(
		a => pp2(2),
		b => pp3(0),
		cin => pp43(4),
		s => pp46(4),
		cout => pp45(5)
		);

	FA421: full_adder port map(
		a => pp2(3),
		b => pp43(5),
		cin => pp44(5),
		s => pp46(5),
		cout => pp45(6)
		);

	FA422: full_adder port map(
		a => pp39(6),
		b => pp43(6),
		cin => pp44(6),
		s => pp46(6),
		cout => pp45(7)
		);

	FA423: full_adder port map(
		a => pp40(7),
		b => pp43(7),
		cin => pp44(7),
		s => pp46(7),
		cout => pp45(8)
		);

	FA424: full_adder port map(
		a => pp41(8),
		b => pp43(8),
		cin => pp44(8),
		s => pp46(8),
		cout => pp45(9)
		);

	FA425: full_adder port map(
		a => pp42(9),
		b => pp43(9),
		cin => pp44(9),
		s => pp46(9),
		cout => pp45(10)
		);

	FA426: full_adder port map(
		a => pp42(10),
		b => pp43(10),
		cin => pp44(10),
		s => pp46(10),
		cout => pp45(11)
		);

	FA427: full_adder port map(
		a => pp42(11),
		b => pp43(11),
		cin => pp44(11),
		s => pp46(11),
		cout => pp45(12)
		);

	FA428: full_adder port map(
		a => pp42(12),
		b => pp43(12),
		cin => pp44(12),
		s => pp46(12),
		cout => pp45(13)
		);

	FA429: full_adder port map(
		a => pp42(13),
		b => pp43(13),
		cin => pp44(13),
		s => pp46(13),
		cout => pp45(14)
		);

	FA430: full_adder port map(
		a => pp42(14),
		b => pp43(14),
		cin => pp44(14),
		s => pp46(14),
		cout => pp45(15)
		);

	FA431: full_adder port map(
		a => pp42(15),
		b => pp43(15),
		cin => pp44(15),
		s => pp46(15),
		cout => pp45(16)
		);

	FA432: full_adder port map(
		a => pp42(16),
		b => pp43(16),
		cin => pp44(16),
		s => pp46(16),
		cout => pp45(17)
		);

	FA433: full_adder port map(
		a => pp42(17),
		b => pp43(17),
		cin => pp44(17),
		s => pp46(17),
		cout => pp45(18)
		);

	FA434: full_adder port map(
		a => pp42(18),
		b => pp43(18),
		cin => pp44(18),
		s => pp46(18),
		cout => pp45(19)
		);

	FA435: full_adder port map(
		a => pp42(19),
		b => pp43(19),
		cin => pp44(19),
		s => pp46(19),
		cout => pp45(20)
		);

	FA436: full_adder port map(
		a => pp42(20),
		b => pp43(20),
		cin => pp44(20),
		s => pp46(20),
		cout => pp45(21)
		);

	FA437: full_adder port map(
		a => pp42(21),
		b => pp43(21),
		cin => pp44(21),
		s => pp46(21),
		cout => pp45(22)
		);

	FA438: full_adder port map(
		a => pp42(22),
		b => pp43(22),
		cin => pp44(22),
		s => pp46(22),
		cout => pp45(23)
		);

	FA439: full_adder port map(
		a => pp42(23),
		b => pp43(23),
		cin => pp44(23),
		s => pp46(23),
		cout => pp45(24)
		);

	FA440: full_adder port map(
		a => pp42(24),
		b => pp43(24),
		cin => pp44(24),
		s => pp46(24),
		cout => pp45(25)
		);

	FA441: full_adder port map(
		a => pp42(25),
		b => pp43(25),
		cin => pp44(25),
		s => pp46(25),
		cout => pp45(26)
		);

	FA442: full_adder port map(
		a => pp42(26),
		b => pp43(26),
		cin => pp44(26),
		s => pp46(26),
		cout => pp45(27)
		);

	FA443: full_adder port map(
		a => pp42(27),
		b => pp43(27),
		cin => pp44(27),
		s => pp46(27),
		cout => pp45(28)
		);

	FA444: full_adder port map(
		a => pp42(28),
		b => pp43(28),
		cin => pp44(28),
		s => pp46(28),
		cout => pp45(29)
		);

	FA445: full_adder port map(
		a => pp42(29),
		b => pp43(29),
		cin => pp44(29),
		s => pp46(29),
		cout => pp45(30)
		);

	FA446: full_adder port map(
		a => pp42(30),
		b => pp43(30),
		cin => pp44(30),
		s => pp46(30),
		cout => pp45(31)
		);

	FA447: full_adder port map(
		a => pp42(31),
		b => pp43(31),
		cin => pp44(31),
		s => pp46(31),
		cout => pp45(32)
		);

	FA448: full_adder port map(
		a => pp42(32),
		b => pp43(32),
		cin => pp44(32),
		s => pp46(32),
		cout => pp45(33)
		);

	FA449: full_adder port map(
		a => pp42(33),
		b => pp43(33),
		cin => pp44(33),
		s => pp46(33),
		cout => pp45(34)
		);

	FA450: full_adder port map(
		a => pp42(34),
		b => pp43(34),
		cin => pp44(34),
		s => pp46(34),
		cout => pp45(35)
		);

	FA451: full_adder port map(
		a => pp42(35),
		b => pp43(35),
		cin => pp44(35),
		s => pp46(35),
		cout => pp45(36)
		);

	FA452: full_adder port map(
		a => pp42(36),
		b => pp43(36),
		cin => pp44(36),
		s => pp46(36),
		cout => pp45(37)
		);

	FA453: full_adder port map(
		a => pp42(37),
		b => pp43(37),
		cin => pp44(37),
		s => pp46(37),
		cout => pp45(38)
		);

	FA454: full_adder port map(
		a => pp42(38),
		b => pp43(38),
		cin => pp44(38),
		s => pp46(38),
		cout => pp45(39)
		);

	FA455: full_adder port map(
		a => pp42(39),
		b => pp43(39),
		cin => pp44(39),
		s => pp46(39),
		cout => pp45(40)
		);

	FA456: full_adder port map(
		a => pp42(40),
		b => pp43(40),
		cin => pp44(40),
		s => pp46(40),
		cout => pp45(41)
		);

	FA457: full_adder port map(
		a => pp42(41),
		b => pp43(41),
		cin => pp44(41),
		s => pp46(41),
		cout => pp45(42)
		);

	FA458: full_adder port map(
		a => pp42(42),
		b => pp43(42),
		cin => pp44(42),
		s => pp46(42),
		cout => pp45(43)
		);

	FA459: full_adder port map(
		a => pp42(43),
		b => pp43(43),
		cin => pp44(43),
		s => pp46(43),
		cout => pp45(44)
		);

	FA460: full_adder port map(
		a => pp42(44),
		b => pp43(44),
		cin => pp44(44),
		s => pp46(44),
		cout => pp45(45)
		);

	FA461: full_adder port map(
		a => pp42(45),
		b => pp43(45),
		cin => pp44(45),
		s => pp46(45),
		cout => pp45(46)
		);

	FA462: full_adder port map(
		a => pp42(46),
		b => pp43(46),
		cin => pp44(46),
		s => pp46(46),
		cout => pp45(47)
		);

	FA463: full_adder port map(
		a => pp42(47),
		b => pp43(47),
		cin => pp44(47),
		s => pp46(47),
		cout => pp45(48)
		);

	FA464: full_adder port map(
		a => pp42(48),
		b => pp43(48),
		cin => pp44(48),
		s => pp46(48),
		cout => pp45(49)
		);

	FA465: full_adder port map(
		a => pp42(49),
		b => pp43(49),
		cin => pp44(49),
		s => pp46(49),
		cout => pp45(50)
		);

	FA466: full_adder port map(
		a => pp42(50),
		b => pp43(50),
		cin => pp44(50),
		s => pp46(50),
		cout => pp45(51)
		);

	FA467: full_adder port map(
		a => pp42(51),
		b => pp43(51),
		cin => pp44(51),
		s => pp46(51),
		cout => pp45(52)
		);

	FA468: full_adder port map(
		a => pp42(52),
		b => pp43(52),
		cin => pp44(52),
		s => pp46(52),
		cout => pp45(53)
		);

	FA469: full_adder port map(
		a => pp42(53),
		b => pp43(53),
		cin => pp44(53),
		s => pp46(53),
		cout => pp45(54)
		);

	FA470: full_adder port map(
		a => pp42(54),
		b => pp43(54),
		cin => pp44(54),
		s => pp46(54),
		cout => pp45(55)
		);

	FA471: full_adder port map(
		a => pp42(55),
		b => pp43(55),
		cin => pp44(55),
		s => pp46(55),
		cout => pp45(56)
		);

	FA472: full_adder port map(
		a => pp42(56),
		b => pp43(56),
		cin => pp44(56),
		s => pp46(56),
		cout => pp45(57)
		);

	FA473: full_adder port map(
		a => pp42(57),
		b => pp43(57),
		cin => pp44(57),
		s => pp46(57),
		cout => pp45(58)
		);

	FA474: full_adder port map(
		a => pp42(58),
		b => pp43(58),
		cin => pp44(58),
		s => pp46(58),
		cout => pp45(59)
		);

	FA475: full_adder port map(
		a => pp41(59),
		b => pp43(59),
		cin => pp44(59),
		s => pp46(59),
		cout => pp45(60)
		);

	FA476: full_adder port map(
		a => pp40(60),
		b => pp43(60),
		cin => pp44(60),
		s => pp46(60),
		cout => pp45(61)
		);

	FA477: full_adder port map(
		a => pp39(61),
		b => pp43(61),
		cin => pp44(61),
		s => pp46(61),
		cout => pp45(62)
		);

	FA478: full_adder port map(
		a => pp16(32),
		b => pp43(62),
		cin => pp44(62),
		s => pp46(62),
		cout => pp45(63)
		);

	FA479: full_adder port map(
		a => pp15(35),
		b => pp16(33),
		cin => pp43(63),
		s => pp46(63),
		cout => open
		);

	pp45(0) <= pp0(0);
	pp45(1) <= pp0(1);
	pp46(0) <= pp1(0);
	pp46(2) <= pp2(0);
	final0(0) <= pp45(0);
	final1(0) <= pp46(0);
	final0(1) <= pp45(1);
	final1(1) <= '0';
	final0(2) <= pp45(2);
	final1(2) <= pp46(2);
	final0(3) <= pp45(3);
	final1(3) <= pp46(3);
	final0(4) <= pp45(4);
	final1(4) <= pp46(4);
	final0(5) <= pp45(5);
	final1(5) <= pp46(5);
	final0(6) <= pp45(6);
	final1(6) <= pp46(6);
	final0(7) <= pp45(7);
	final1(7) <= pp46(7);
	final0(8) <= pp45(8);
	final1(8) <= pp46(8);
	final0(9) <= pp45(9);
	final1(9) <= pp46(9);
	final0(10) <= pp45(10);
	final1(10) <= pp46(10);
	final0(11) <= pp45(11);
	final1(11) <= pp46(11);
	final0(12) <= pp45(12);
	final1(12) <= pp46(12);
	final0(13) <= pp45(13);
	final1(13) <= pp46(13);
	final0(14) <= pp45(14);
	final1(14) <= pp46(14);
	final0(15) <= pp45(15);
	final1(15) <= pp46(15);
	final0(16) <= pp45(16);
	final1(16) <= pp46(16);
	final0(17) <= pp45(17);
	final1(17) <= pp46(17);
	final0(18) <= pp45(18);
	final1(18) <= pp46(18);
	final0(19) <= pp45(19);
	final1(19) <= pp46(19);
	final0(20) <= pp45(20);
	final1(20) <= pp46(20);
	final0(21) <= pp45(21);
	final1(21) <= pp46(21);
	final0(22) <= pp45(22);
	final1(22) <= pp46(22);
	final0(23) <= pp45(23);
	final1(23) <= pp46(23);
	final0(24) <= pp45(24);
	final1(24) <= pp46(24);
	final0(25) <= pp45(25);
	final1(25) <= pp46(25);
	final0(26) <= pp45(26);
	final1(26) <= pp46(26);
	final0(27) <= pp45(27);
	final1(27) <= pp46(27);
	final0(28) <= pp45(28);
	final1(28) <= pp46(28);
	final0(29) <= pp45(29);
	final1(29) <= pp46(29);
	final0(30) <= pp45(30);
	final1(30) <= pp46(30);
	final0(31) <= pp45(31);
	final1(31) <= pp46(31);
	final0(32) <= pp45(32);
	final1(32) <= pp46(32);
	final0(33) <= pp45(33);
	final1(33) <= pp46(33);
	final0(34) <= pp45(34);
	final1(34) <= pp46(34);
	final0(35) <= pp45(35);
	final1(35) <= pp46(35);
	final0(36) <= pp45(36);
	final1(36) <= pp46(36);
	final0(37) <= pp45(37);
	final1(37) <= pp46(37);
	final0(38) <= pp45(38);
	final1(38) <= pp46(38);
	final0(39) <= pp45(39);
	final1(39) <= pp46(39);
	final0(40) <= pp45(40);
	final1(40) <= pp46(40);
	final0(41) <= pp45(41);
	final1(41) <= pp46(41);
	final0(42) <= pp45(42);
	final1(42) <= pp46(42);
	final0(43) <= pp45(43);
	final1(43) <= pp46(43);
	final0(44) <= pp45(44);
	final1(44) <= pp46(44);
	final0(45) <= pp45(45);
	final1(45) <= pp46(45);
	final0(46) <= pp45(46);
	final1(46) <= pp46(46);
	final0(47) <= pp45(47);
	final1(47) <= pp46(47);
	final0(48) <= pp45(48);
	final1(48) <= pp46(48);
	final0(49) <= pp45(49);
	final1(49) <= pp46(49);
	final0(50) <= pp45(50);
	final1(50) <= pp46(50);
	final0(51) <= pp45(51);
	final1(51) <= pp46(51);
	final0(52) <= pp45(52);
	final1(52) <= pp46(52);
	final0(53) <= pp45(53);
	final1(53) <= pp46(53);
	final0(54) <= pp45(54);
	final1(54) <= pp46(54);
	final0(55) <= pp45(55);
	final1(55) <= pp46(55);
	final0(56) <= pp45(56);
	final1(56) <= pp46(56);
	final0(57) <= pp45(57);
	final1(57) <= pp46(57);
	final0(58) <= pp45(58);
	final1(58) <= pp46(58);
	final0(59) <= pp45(59);
	final1(59) <= pp46(59);
	final0(60) <= pp45(60);
	final1(60) <= pp46(60);
	final0(61) <= pp45(61);
	final1(61) <= pp46(61);
	final0(62) <= pp45(62);
	final1(62) <= pp46(62);
	final0(63) <= pp45(63);
	final1(63) <= pp46(63);

end structural;
