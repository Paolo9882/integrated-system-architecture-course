library verilog;
use verilog.vl_types.all;
entity tb_FPmul is
end tb_FPmul;
